// Verilog netlist created by TD v5.0.31956
// Wed Dec  1 01:17:01 2021

`timescale 1ns / 1ps
module rom0  // rom0.v(14)
  (
  addra,
  clka,
  rsta,
  doa
  );

  input [12:0] addra;  // rom0.v(18)
  input clka;  // rom0.v(19)
  input rsta;  // rom0.v(20)
  output [31:0] doa;  // rom0.v(16)

  wire [0:2] addra_piped;
  wire  \inst_doa_mux_b0/B0_0 ;
  wire  \inst_doa_mux_b0/B0_1 ;
  wire  \inst_doa_mux_b0/B0_2 ;
  wire  \inst_doa_mux_b0/B0_3 ;
  wire  \inst_doa_mux_b0/B1_0 ;
  wire  \inst_doa_mux_b0/B1_1 ;
  wire  \inst_doa_mux_b1/B0_0 ;
  wire  \inst_doa_mux_b1/B0_1 ;
  wire  \inst_doa_mux_b1/B0_2 ;
  wire  \inst_doa_mux_b1/B0_3 ;
  wire  \inst_doa_mux_b1/B1_0 ;
  wire  \inst_doa_mux_b1/B1_1 ;
  wire  \inst_doa_mux_b10/B0_0 ;
  wire  \inst_doa_mux_b10/B1_0 ;
  wire  \inst_doa_mux_b11/B0_0 ;
  wire  \inst_doa_mux_b11/B0_1 ;
  wire  \inst_doa_mux_b11/B0_2 ;
  wire  \inst_doa_mux_b11/B0_3 ;
  wire  \inst_doa_mux_b11/B1_0 ;
  wire  \inst_doa_mux_b11/B1_1 ;
  wire  \inst_doa_mux_b12/B0_0 ;
  wire  \inst_doa_mux_b12/B0_1 ;
  wire  \inst_doa_mux_b12/B0_2 ;
  wire  \inst_doa_mux_b12/B0_3 ;
  wire  \inst_doa_mux_b12/B1_0 ;
  wire  \inst_doa_mux_b12/B1_1 ;
  wire  \inst_doa_mux_b13/B0_0 ;
  wire  \inst_doa_mux_b13/B0_1 ;
  wire  \inst_doa_mux_b13/B0_2 ;
  wire  \inst_doa_mux_b13/B0_3 ;
  wire  \inst_doa_mux_b13/B1_0 ;
  wire  \inst_doa_mux_b13/B1_1 ;
  wire  \inst_doa_mux_b14/B0_0 ;
  wire  \inst_doa_mux_b14/B0_1 ;
  wire  \inst_doa_mux_b14/B0_2 ;
  wire  \inst_doa_mux_b14/B0_3 ;
  wire  \inst_doa_mux_b14/B1_0 ;
  wire  \inst_doa_mux_b14/B1_1 ;
  wire  \inst_doa_mux_b15/B0_0 ;
  wire  \inst_doa_mux_b15/B0_1 ;
  wire  \inst_doa_mux_b15/B0_2 ;
  wire  \inst_doa_mux_b15/B0_3 ;
  wire  \inst_doa_mux_b15/B1_0 ;
  wire  \inst_doa_mux_b15/B1_1 ;
  wire  \inst_doa_mux_b16/B0_0 ;
  wire  \inst_doa_mux_b16/B0_1 ;
  wire  \inst_doa_mux_b16/B0_2 ;
  wire  \inst_doa_mux_b16/B0_3 ;
  wire  \inst_doa_mux_b16/B1_0 ;
  wire  \inst_doa_mux_b16/B1_1 ;
  wire  \inst_doa_mux_b17/B0_0 ;
  wire  \inst_doa_mux_b17/B0_1 ;
  wire  \inst_doa_mux_b17/B0_2 ;
  wire  \inst_doa_mux_b17/B0_3 ;
  wire  \inst_doa_mux_b17/B1_0 ;
  wire  \inst_doa_mux_b17/B1_1 ;
  wire  \inst_doa_mux_b18/B0_0 ;
  wire  \inst_doa_mux_b18/B1_0 ;
  wire  \inst_doa_mux_b2/B0_0 ;
  wire  \inst_doa_mux_b2/B1_0 ;
  wire  \inst_doa_mux_b3/B0_0 ;
  wire  \inst_doa_mux_b3/B1_0 ;
  wire  \inst_doa_mux_b4/B0_0 ;
  wire  \inst_doa_mux_b4/B1_0 ;
  wire  \inst_doa_mux_b5/B0_0 ;
  wire  \inst_doa_mux_b5/B1_0 ;
  wire  \inst_doa_mux_b6/B0_0 ;
  wire  \inst_doa_mux_b6/B1_0 ;
  wire  \inst_doa_mux_b7/B0_0 ;
  wire  \inst_doa_mux_b7/B1_0 ;
  wire  \inst_doa_mux_b8/B0_0 ;
  wire  \inst_doa_mux_b8/B1_0 ;
  wire inst_doa_i0_000;
  wire inst_doa_i0_001;
  wire inst_doa_i0_002;
  wire inst_doa_i0_003;
  wire inst_doa_i0_004;
  wire inst_doa_i0_005;
  wire inst_doa_i0_006;
  wire inst_doa_i0_007;
  wire inst_doa_i0_008;
  wire inst_doa_i0_009;
  wire inst_doa_i0_010;
  wire inst_doa_i0_011;
  wire inst_doa_i0_012;
  wire inst_doa_i0_013;
  wire inst_doa_i0_014;
  wire inst_doa_i0_015;
  wire inst_doa_i0_016;
  wire inst_doa_i0_017;
  wire inst_doa_i0_027;
  wire inst_doa_i1_000;
  wire inst_doa_i1_001;
  wire inst_doa_i1_002;
  wire inst_doa_i1_003;
  wire inst_doa_i1_004;
  wire inst_doa_i1_005;
  wire inst_doa_i1_006;
  wire inst_doa_i1_007;
  wire inst_doa_i1_008;
  wire inst_doa_i2_000;
  wire inst_doa_i2_001;
  wire inst_doa_i2_002;
  wire inst_doa_i2_003;
  wire inst_doa_i2_004;
  wire inst_doa_i2_005;
  wire inst_doa_i2_006;
  wire inst_doa_i2_007;
  wire inst_doa_i2_008;
  wire inst_doa_i3_000;
  wire inst_doa_i3_001;
  wire inst_doa_i3_002;
  wire inst_doa_i3_003;
  wire inst_doa_i3_004;
  wire inst_doa_i3_005;
  wire inst_doa_i3_006;
  wire inst_doa_i3_007;
  wire inst_doa_i3_008;
  wire inst_doa_i4_000;
  wire inst_doa_i4_001;
  wire inst_doa_i4_002;
  wire inst_doa_i4_003;
  wire inst_doa_i4_004;
  wire inst_doa_i4_005;
  wire inst_doa_i4_006;
  wire inst_doa_i4_007;
  wire inst_doa_i4_008;
  wire inst_doa_i5_000;
  wire inst_doa_i5_001;
  wire inst_doa_i5_002;
  wire inst_doa_i5_003;
  wire inst_doa_i5_004;
  wire inst_doa_i5_005;
  wire inst_doa_i5_006;
  wire inst_doa_i5_007;
  wire inst_doa_i5_008;
  wire inst_doa_i6_000;
  wire inst_doa_i6_001;
  wire inst_doa_i6_002;
  wire inst_doa_i6_003;
  wire inst_doa_i6_004;
  wire inst_doa_i6_005;
  wire inst_doa_i6_006;
  wire inst_doa_i6_007;
  wire inst_doa_i6_008;
  wire inst_doa_i7_000;
  wire inst_doa_i7_001;
  wire inst_doa_i7_002;
  wire inst_doa_i7_003;
  wire inst_doa_i7_004;
  wire inst_doa_i7_005;
  wire inst_doa_i7_006;
  wire inst_doa_i7_007;
  wire inst_doa_i7_008;

  assign doa[31] = inst_doa_i0_027;
  assign doa[30] = inst_doa_i0_027;
  assign doa[29] = inst_doa_i0_027;
  assign doa[28] = inst_doa_i0_027;
  assign doa[27] = inst_doa_i0_027;
  assign doa[26] = doa[17];
  assign doa[25] = doa[16];
  assign doa[24] = doa[15];
  assign doa[23] = doa[14];
  assign doa[22] = doa[13];
  assign doa[21] = doa[12];
  assign doa[20] = doa[11];
  assign doa[19] = doa[10];
  assign doa[9] = doa[18];
  AL_DFF_X addra_pipe_b0 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clka),
    .d(addra[10]),
    .en(1'b1),
    .sr(rsta),
    .ss(1'b0),
    .q(addra_piped[0]));
  AL_DFF_X addra_pipe_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clka),
    .d(addra[11]),
    .en(1'b1),
    .sr(rsta),
    .ss(1'b0),
    .q(addra_piped[1]));
  AL_DFF_X addra_pipe_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clka),
    .d(addra[12]),
    .en(1'b1),
    .sr(rsta),
    .ss(1'b0),
    .q(addra_piped[2]));
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h000000000000000000000000000000000000008067130313132313676F6F6F37),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i0_008,inst_doa_i0_007,inst_doa_i0_006,inst_doa_i0_005,inst_doa_i0_004,inst_doa_i0_003,inst_doa_i0_002,inst_doa_i0_001,inst_doa_i0_000}));
  // address_offset=0;data_offset=9;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_009 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i0_017,inst_doa_i0_016,inst_doa_i0_015,inst_doa_i0_014,inst_doa_i0_013,inst_doa_i0_012,inst_doa_i0_011,inst_doa_i0_010,inst_doa_i0_009}));
  // address_offset=0;data_offset=27;depth=8192;width=1;num_section=1;width_per_section=1;section_size=32;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("1"),
    .CSA1("1"),
    .CSA2("1"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_000000_027 (
    .addra(addra),
    .clka(clka),
    .dia({open_n153,open_n154,open_n155,open_n156,open_n157,open_n158,open_n159,1'b0,open_n160}),
    .rsta(rsta),
    .doa({open_n175,open_n176,open_n177,open_n178,open_n179,open_n180,open_n181,open_n182,inst_doa_i0_027}));
  // address_offset=1024;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_001024_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i1_008,inst_doa_i1_007,inst_doa_i1_006,inst_doa_i1_005,inst_doa_i1_004,inst_doa_i1_003,inst_doa_i1_002,inst_doa_i1_001,inst_doa_i1_000}));
  // address_offset=2048;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_002048_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i2_008,inst_doa_i2_007,inst_doa_i2_006,inst_doa_i2_005,inst_doa_i2_004,inst_doa_i2_003,inst_doa_i2_002,inst_doa_i2_001,inst_doa_i2_000}));
  // address_offset=3072;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_003072_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i3_008,inst_doa_i3_007,inst_doa_i3_006,inst_doa_i3_005,inst_doa_i3_004,inst_doa_i3_003,inst_doa_i3_002,inst_doa_i3_001,inst_doa_i3_000}));
  // address_offset=4096;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_004096_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i4_008,inst_doa_i4_007,inst_doa_i4_006,inst_doa_i4_005,inst_doa_i4_004,inst_doa_i4_003,inst_doa_i4_002,inst_doa_i4_001,inst_doa_i4_000}));
  // address_offset=5120;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_005120_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i5_008,inst_doa_i5_007,inst_doa_i5_006,inst_doa_i5_005,inst_doa_i5_004,inst_doa_i5_003,inst_doa_i5_002,inst_doa_i5_001,inst_doa_i5_000}));
  // address_offset=6144;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_006144_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i6_008,inst_doa_i6_007,inst_doa_i6_006,inst_doa_i6_005,inst_doa_i6_004,inst_doa_i6_003,inst_doa_i6_002,inst_doa_i6_001,inst_doa_i6_000}));
  // address_offset=7168;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=32;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("0"),
    .CLKBMUX("0"),
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("1"),
    .CSB1("1"),
    .CSB2("1"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .MODE("SP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTBMUX("0"),
    .WEAMUX("0"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_8192x32_sub_007168_000 (
    .addra({addra[9:0],3'b111}),
    .clka(clka),
    .csa(addra[12:10]),
    .dia(9'b000000000),
    .rsta(rsta),
    .doa({inst_doa_i7_008,inst_doa_i7_007,inst_doa_i7_006,inst_doa_i7_005,inst_doa_i7_004,inst_doa_i7_003,inst_doa_i7_002,inst_doa_i7_001,inst_doa_i7_000}));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_0  (
    .i0(inst_doa_i0_000),
    .i1(inst_doa_i1_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_0 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_1  (
    .i0(inst_doa_i2_000),
    .i1(inst_doa_i3_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_1 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_2  (
    .i0(inst_doa_i4_000),
    .i1(inst_doa_i5_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_2 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_0_3  (
    .i0(inst_doa_i6_000),
    .i1(inst_doa_i7_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b0/B0_3 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b0/B0_0 ),
    .i1(\inst_doa_mux_b0/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_0 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b0/B0_2 ),
    .i1(\inst_doa_mux_b0/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b0/B1_1 ));
  AL_MUX \inst_doa_mux_b0/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b0/B1_0 ),
    .i1(\inst_doa_mux_b0/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[0]));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_0  (
    .i0(inst_doa_i0_001),
    .i1(inst_doa_i1_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_0 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_1  (
    .i0(inst_doa_i2_001),
    .i1(inst_doa_i3_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_1 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_2  (
    .i0(inst_doa_i4_001),
    .i1(inst_doa_i5_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_2 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_0_3  (
    .i0(inst_doa_i6_001),
    .i1(inst_doa_i7_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b1/B0_3 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b1/B0_0 ),
    .i1(\inst_doa_mux_b1/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_0 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b1/B0_2 ),
    .i1(\inst_doa_mux_b1/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b1/B1_1 ));
  AL_MUX \inst_doa_mux_b1/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b1/B1_0 ),
    .i1(\inst_doa_mux_b1/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[1]));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_0_0  (
    .i0(inst_doa_i0_010),
    .i1(inst_doa_i1_001),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b10/B0_0 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b10/B0_0 ),
    .i1(\inst_doa_mux_b1/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b10/B1_0 ));
  AL_MUX \inst_doa_mux_b10/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b10/B1_0 ),
    .i1(\inst_doa_mux_b1/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[10]));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_0_0  (
    .i0(inst_doa_i0_011),
    .i1(inst_doa_i1_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b11/B0_0 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_0_1  (
    .i0(inst_doa_i2_002),
    .i1(inst_doa_i3_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b11/B0_1 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_0_2  (
    .i0(inst_doa_i4_002),
    .i1(inst_doa_i5_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b11/B0_2 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_0_3  (
    .i0(inst_doa_i6_002),
    .i1(inst_doa_i7_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b11/B0_3 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b11/B0_0 ),
    .i1(\inst_doa_mux_b11/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b11/B1_0 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b11/B0_2 ),
    .i1(\inst_doa_mux_b11/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b11/B1_1 ));
  AL_MUX \inst_doa_mux_b11/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b11/B1_0 ),
    .i1(\inst_doa_mux_b11/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[11]));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_0_0  (
    .i0(inst_doa_i0_012),
    .i1(inst_doa_i1_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b12/B0_0 ));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_0_1  (
    .i0(inst_doa_i2_003),
    .i1(inst_doa_i3_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b12/B0_1 ));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_0_2  (
    .i0(inst_doa_i4_003),
    .i1(inst_doa_i5_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b12/B0_2 ));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_0_3  (
    .i0(inst_doa_i6_003),
    .i1(inst_doa_i7_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b12/B0_3 ));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b12/B0_0 ),
    .i1(\inst_doa_mux_b12/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b12/B1_0 ));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b12/B0_2 ),
    .i1(\inst_doa_mux_b12/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b12/B1_1 ));
  AL_MUX \inst_doa_mux_b12/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b12/B1_0 ),
    .i1(\inst_doa_mux_b12/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[12]));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_0_0  (
    .i0(inst_doa_i0_013),
    .i1(inst_doa_i1_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b13/B0_0 ));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_0_1  (
    .i0(inst_doa_i2_004),
    .i1(inst_doa_i3_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b13/B0_1 ));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_0_2  (
    .i0(inst_doa_i4_004),
    .i1(inst_doa_i5_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b13/B0_2 ));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_0_3  (
    .i0(inst_doa_i6_004),
    .i1(inst_doa_i7_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b13/B0_3 ));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b13/B0_0 ),
    .i1(\inst_doa_mux_b13/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b13/B1_0 ));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b13/B0_2 ),
    .i1(\inst_doa_mux_b13/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b13/B1_1 ));
  AL_MUX \inst_doa_mux_b13/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b13/B1_0 ),
    .i1(\inst_doa_mux_b13/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[13]));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_0_0  (
    .i0(inst_doa_i0_014),
    .i1(inst_doa_i1_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b14/B0_0 ));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_0_1  (
    .i0(inst_doa_i2_005),
    .i1(inst_doa_i3_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b14/B0_1 ));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_0_2  (
    .i0(inst_doa_i4_005),
    .i1(inst_doa_i5_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b14/B0_2 ));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_0_3  (
    .i0(inst_doa_i6_005),
    .i1(inst_doa_i7_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b14/B0_3 ));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b14/B0_0 ),
    .i1(\inst_doa_mux_b14/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b14/B1_0 ));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b14/B0_2 ),
    .i1(\inst_doa_mux_b14/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b14/B1_1 ));
  AL_MUX \inst_doa_mux_b14/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b14/B1_0 ),
    .i1(\inst_doa_mux_b14/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[14]));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_0_0  (
    .i0(inst_doa_i0_015),
    .i1(inst_doa_i1_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b15/B0_0 ));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_0_1  (
    .i0(inst_doa_i2_006),
    .i1(inst_doa_i3_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b15/B0_1 ));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_0_2  (
    .i0(inst_doa_i4_006),
    .i1(inst_doa_i5_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b15/B0_2 ));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_0_3  (
    .i0(inst_doa_i6_006),
    .i1(inst_doa_i7_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b15/B0_3 ));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b15/B0_0 ),
    .i1(\inst_doa_mux_b15/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b15/B1_0 ));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b15/B0_2 ),
    .i1(\inst_doa_mux_b15/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b15/B1_1 ));
  AL_MUX \inst_doa_mux_b15/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b15/B1_0 ),
    .i1(\inst_doa_mux_b15/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[15]));
  AL_MUX \inst_doa_mux_b16/al_mux_b0_0_0  (
    .i0(inst_doa_i0_016),
    .i1(inst_doa_i1_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b16/B0_0 ));
  AL_MUX \inst_doa_mux_b16/al_mux_b0_0_1  (
    .i0(inst_doa_i2_007),
    .i1(inst_doa_i3_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b16/B0_1 ));
  AL_MUX \inst_doa_mux_b16/al_mux_b0_0_2  (
    .i0(inst_doa_i4_007),
    .i1(inst_doa_i5_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b16/B0_2 ));
  AL_MUX \inst_doa_mux_b16/al_mux_b0_0_3  (
    .i0(inst_doa_i6_007),
    .i1(inst_doa_i7_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b16/B0_3 ));
  AL_MUX \inst_doa_mux_b16/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b16/B0_0 ),
    .i1(\inst_doa_mux_b16/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b16/B1_0 ));
  AL_MUX \inst_doa_mux_b16/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b16/B0_2 ),
    .i1(\inst_doa_mux_b16/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b16/B1_1 ));
  AL_MUX \inst_doa_mux_b16/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b16/B1_0 ),
    .i1(\inst_doa_mux_b16/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[16]));
  AL_MUX \inst_doa_mux_b17/al_mux_b0_0_0  (
    .i0(inst_doa_i0_017),
    .i1(inst_doa_i1_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b17/B0_0 ));
  AL_MUX \inst_doa_mux_b17/al_mux_b0_0_1  (
    .i0(inst_doa_i2_008),
    .i1(inst_doa_i3_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b17/B0_1 ));
  AL_MUX \inst_doa_mux_b17/al_mux_b0_0_2  (
    .i0(inst_doa_i4_008),
    .i1(inst_doa_i5_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b17/B0_2 ));
  AL_MUX \inst_doa_mux_b17/al_mux_b0_0_3  (
    .i0(inst_doa_i6_008),
    .i1(inst_doa_i7_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b17/B0_3 ));
  AL_MUX \inst_doa_mux_b17/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b17/B0_0 ),
    .i1(\inst_doa_mux_b17/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b17/B1_0 ));
  AL_MUX \inst_doa_mux_b17/al_mux_b0_1_1  (
    .i0(\inst_doa_mux_b17/B0_2 ),
    .i1(\inst_doa_mux_b17/B0_3 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b17/B1_1 ));
  AL_MUX \inst_doa_mux_b17/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b17/B1_0 ),
    .i1(\inst_doa_mux_b17/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[17]));
  AL_MUX \inst_doa_mux_b18/al_mux_b0_0_0  (
    .i0(inst_doa_i0_009),
    .i1(inst_doa_i1_000),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b18/B0_0 ));
  AL_MUX \inst_doa_mux_b18/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b18/B0_0 ),
    .i1(\inst_doa_mux_b0/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b18/B1_0 ));
  AL_MUX \inst_doa_mux_b18/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b18/B1_0 ),
    .i1(\inst_doa_mux_b0/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[18]));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_0_0  (
    .i0(inst_doa_i0_002),
    .i1(inst_doa_i1_002),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b2/B0_0 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b2/B0_0 ),
    .i1(\inst_doa_mux_b11/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b2/B1_0 ));
  AL_MUX \inst_doa_mux_b2/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b2/B1_0 ),
    .i1(\inst_doa_mux_b11/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[2]));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_0_0  (
    .i0(inst_doa_i0_003),
    .i1(inst_doa_i1_003),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b3/B0_0 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b3/B0_0 ),
    .i1(\inst_doa_mux_b12/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b3/B1_0 ));
  AL_MUX \inst_doa_mux_b3/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b3/B1_0 ),
    .i1(\inst_doa_mux_b12/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[3]));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_0_0  (
    .i0(inst_doa_i0_004),
    .i1(inst_doa_i1_004),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b4/B0_0 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b4/B0_0 ),
    .i1(\inst_doa_mux_b13/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b4/B1_0 ));
  AL_MUX \inst_doa_mux_b4/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b4/B1_0 ),
    .i1(\inst_doa_mux_b13/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[4]));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_0_0  (
    .i0(inst_doa_i0_005),
    .i1(inst_doa_i1_005),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b5/B0_0 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b5/B0_0 ),
    .i1(\inst_doa_mux_b14/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b5/B1_0 ));
  AL_MUX \inst_doa_mux_b5/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b5/B1_0 ),
    .i1(\inst_doa_mux_b14/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[5]));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_0_0  (
    .i0(inst_doa_i0_006),
    .i1(inst_doa_i1_006),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b6/B0_0 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b6/B0_0 ),
    .i1(\inst_doa_mux_b15/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b6/B1_0 ));
  AL_MUX \inst_doa_mux_b6/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b6/B1_0 ),
    .i1(\inst_doa_mux_b15/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[6]));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_0_0  (
    .i0(inst_doa_i0_007),
    .i1(inst_doa_i1_007),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b7/B0_0 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b7/B0_0 ),
    .i1(\inst_doa_mux_b16/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b7/B1_0 ));
  AL_MUX \inst_doa_mux_b7/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b7/B1_0 ),
    .i1(\inst_doa_mux_b16/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[7]));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_0_0  (
    .i0(inst_doa_i0_008),
    .i1(inst_doa_i1_008),
    .sel(addra_piped[0]),
    .o(\inst_doa_mux_b8/B0_0 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_1_0  (
    .i0(\inst_doa_mux_b8/B0_0 ),
    .i1(\inst_doa_mux_b17/B0_1 ),
    .sel(addra_piped[1]),
    .o(\inst_doa_mux_b8/B1_0 ));
  AL_MUX \inst_doa_mux_b8/al_mux_b0_2_0  (
    .i0(\inst_doa_mux_b8/B1_0 ),
    .i1(\inst_doa_mux_b17/B1_1 ),
    .sel(addra_piped[2]),
    .o(doa[8]));

endmodule 

module AL_DFF_X
  (
  ar,
  as,
  clk,
  d,
  en,
  sr,
  ss,
  q
  );

  input ar;
  input as;
  input clk;
  input d;
  input en;
  input sr;
  input ss;
  output q;

  wire enout;
  wire srout;
  wire ssout;

  AL_MUX u_en (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset (
    .i0(ssout),
    .i1(1'b0),
    .sel(sr),
    .o(srout));
  AL_DFF u_seq (
    .clk(clk),
    .d(srout),
    .reset(ar),
    .set(as),
    .q(q));
  AL_MUX u_set (
    .i0(enout),
    .i1(1'b1),
    .sel(ss),
    .o(ssout));

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  // synthesis translate_off
  tri0 gsrn = glbl.gsrn;

  always @(gsrn)
  begin
    if(!gsrn)
      assign q = INI;
    else
      deassign q;
  end
  // synthesis translate_on

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

